library verilog;
use verilog.vl_types.all;
entity tb_inst_mem is
end tb_inst_mem;
