library verilog;
use verilog.vl_types.all;
entity tb_mips is
end tb_mips;
